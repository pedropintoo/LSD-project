library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity NoisyTriangSignal_ROM_256x8 is
   port(address : in  std_logic_vector(7 downto 0);
        dataOut : out std_logic_vector(7 downto 0));
end NoisyTriangSignal_ROM_256x8;

architecture Behavioral of NoisyTriangSignal_ROM_256x8 is
   subtype TDataWord is std_logic_vector(7 downto 0);
   type TROM is array (0 to 255) of TDataWord;
	-- Input Signal ROM
   constant c_memory: TROM := (
		"10110011", -- -77
		"10001110", -- -114
		"10111100", -- -68
		"10101101", -- -83
		"10110110", -- -74
		"10100000", -- -96
		"10101110", -- -82
		"10110100", -- -76
		"10111110", -- -66
		"10101101", -- -83
		"11000101", -- -59
		"10111000", -- -72
		"11000111", -- -57
		"11010000", -- -48
		"11010000", -- -48
		"11011010", -- -38
		"11011101", -- -35
		"11010000", -- -48
		"11011100", -- -36
		"11010100", -- -44
		"11010011", -- -45
		"11101100", -- -20
		"11100110", -- -26
		"11101001", -- -23
		"11110110", -- -10
		"11110110", -- -10
		"11110111", -- -9
		"00000010", -- 2
		"00000011", -- 3
		"11111111", -- -1
		"11111001", -- -7
		"11111101", -- -3
		"00010010", -- 18
		"11111010", -- -6
		"00001101", -- 13
		"11111101", -- -3
		"00011101", -- 29
		"00011111", -- 31
		"00011010", -- 26
		"00011100", -- 28
		"00001000", -- 8
		"00101001", -- 41
		"00010001", -- 17
		"00010011", -- 19
		"00101110", -- 46
		"00100111", -- 39
		"00110111", -- 55
		"00111101", -- 61
		"01000010", -- 66
		"00110110", -- 54
		"01000100", -- 68
		"01000100", -- 68
		"01001110", -- 78
		"01001111", -- 79
		"01010101", -- 85
		"01001111", -- 79
		"01010010", -- 82
		"01100000", -- 96
		"01000101", -- 69
		"01011000", -- 88
		"01010100", -- 84
		"01011001", -- 89
		"01100000", -- 96
		"01011110", -- 94
		"01001001", -- 73
		"01001011", -- 75
		"01001110", -- 78
		"01000111", -- 71
		"01001001", -- 73
		"01000111", -- 71
		"00110111", -- 55
		"00111011", -- 59
		"00100101", -- 37
		"01000001", -- 65
		"00101101", -- 45
		"00100100", -- 36
		"00101010", -- 42
		"00011100", -- 28
		"00100110", -- 38
		"00011110", -- 30
		"00110101", -- 53
		"00101000", -- 40
		"00000010", -- 2
		"00011011", -- 27
		"00000110", -- 6
		"00001110", -- 14
		"00001110", -- 14
		"00010001", -- 17
		"00000100", -- 4
		"00010010", -- 18
		"11111011", -- -5
		"00000000", -- 0
		"00000000", -- 0
		"11110111", -- -9
		"11111100", -- -4
		"11110011", -- -13
		"11100101", -- -27
		"11011000", -- -40
		"11111000", -- -8
		"11011101", -- -35
		"11100001", -- -31
		"11100010", -- -30
		"11011011", -- -37
		"11001110", -- -50
		"11001111", -- -49
		"11001111", -- -49
		"11011011", -- -37
		"11000001", -- -63
		"11001110", -- -50
		"11000110", -- -58
		"10111110", -- -66
		"10110011", -- -77
		"10110111", -- -73
		"10110110", -- -74
		"10100101", -- -91
		"10110010", -- -78
		"10100101", -- -91
		"10101001", -- -87
		"10101010", -- -86
		"10011011", -- -101
		"10011101", -- -99
		"10100111", -- -89
		"10010101", -- -107
		"10110100", -- -76
		"11000100", -- -60
		"10111001", -- -71
		"10110000", -- -80
		"10111011", -- -69
		"10110000", -- -80
		"11001111", -- -49
		"11001001", -- -55
		"11001011", -- -53
		"10111110", -- -66
		"11001101", -- -51
		"11000111", -- -57
		"11001101", -- -51
		"11001110", -- -50
		"11001101", -- -51
		"11010001", -- -47
		"11011011", -- -37
		"11010000", -- -48
		"11101001", -- -23
		"11100101", -- -27
		"11110000", -- -16
		"11101111", -- -17
		"11110101", -- -11
		"11100101", -- -27
		"11101101", -- -19
		"11110101", -- -11
		"11111110", -- -2
		"00001011", -- 11
		"00000000", -- 0
		"00010011", -- 19
		"00001110", -- 14
		"00011000", -- 24
		"00010001", -- 17
		"00001101", -- 13
		"00001000", -- 8
		"00011011", -- 27
		"00100101", -- 37
		"00011101", -- 29
		"00011110", -- 30
		"00100011", -- 35
		"00011111", -- 31
		"00101000", -- 40
		"00101110", -- 46
		"00110100", -- 52
		"00110110", -- 54
		"00111111", -- 63
		"00111110", -- 62
		"01010001", -- 81
		"01000110", -- 70
		"01011000", -- 88
		"01000011", -- 67
		"01010010", -- 82
		"01001110", -- 78
		"01011001", -- 89
		"01011100", -- 92
		"01000101", -- 69
		"01010000", -- 80
		"01010010", -- 82
		"01100001", -- 97
		"01101000", -- 104
		"01010011", -- 83
		"01011011", -- 91
		"01010101", -- 85
		"01000011", -- 67
		"01001101", -- 77
		"00111111", -- 63
		"01010010", -- 82
		"01000000", -- 64
		"01001101", -- 77
		"00110110", -- 54
		"00111100", -- 60
		"00110011", -- 51
		"00011101", -- 29
		"00100011", -- 35
		"00101111", -- 47
		"00100110", -- 38
		"00011000", -- 24
		"00011010", -- 26
		"00011111", -- 31
		"00010000", -- 16
		"00100000", -- 32
		"00001101", -- 13
		"00100001", -- 33
		"00000010", -- 2
		"00001100", -- 12
		"11111000", -- -8
		"11111100", -- -4
		"11111010", -- -6
		"00000001", -- 1
		"00000011", -- 3
		"11111001", -- -7
		"11110000", -- -16
		"11111000", -- -8
		"11110100", -- -12
		"11101011", -- -21
		"11101100", -- -20
		"11100111", -- -25
		"11010111", -- -41
		"11100100", -- -28
		"11010011", -- -45
		"11010001", -- -47
		"11010101", -- -43
		"11001101", -- -51
		"11001100", -- -52
		"11001111", -- -49
		"11010000", -- -48
		"11000001", -- -63
		"11000011", -- -61
		"10111011", -- -69
		"10111100", -- -68
		"10111011", -- -69
		"10101101", -- -83
		"10110011", -- -77
		"10110011", -- -77
		"10101010", -- -86
		"10110111", -- -73
		"10011101", -- -99
		"10011001", -- -103
		"10010010", -- -110
		"10101111", -- -81
		"10110010", -- -78
		"10101100", -- -84
		"10111001", -- -71
		"10110101", -- -75
		"10111001", -- -71
		"10111011", -- -69
		"11000001", -- -63
		"11000001", -- -63
		"11011110", -- -34
		"10111011", -- -69
		"10111000", -- -72
		"11000010", -- -62
		"11000110" -- -58
);

begin
   dataOut <= c_memory(to_integer(unsigned(address)));
end Behavioral;
